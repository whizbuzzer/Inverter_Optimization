A simple AC run - this is just a comment!
.options list node post
.op
.ac dec 10 1k 1x
.print ac v(1) v(2) i(r2) i(c1)
v1 1 0 10 ac 1
r1 1 2 1k
r2 2 0 1k
c1 2 0 .001u
.end
